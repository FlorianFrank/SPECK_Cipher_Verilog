`ifndef _general_settings_
`define _general_settings_

	//% Number of rounds to be executed.
	`define NR_ROUNDS 32'd31
	//% The key size in bits.
	`define KEY_SIZE 32'd128
	//% The block size in bits.
	`define BLOCK_SIZE 32'd64

`endif //_general_settings_
