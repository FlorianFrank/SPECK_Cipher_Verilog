`ifndef _main_module_defines_
`define _main_module_defines_

`define WAIT_FOR_START_SIGNAL 	        0
`define START_KEY_SCHEDULE  		    1
`define STOP_KEY_SCHEDULE 			    2
`define START_ROUND  				    3
`define STOP_ROUND 					    4
`define ITERATE_CTR 					5
`define DONE 							6

`define CACHE_ROUND_KEYS                7
`endif // _main_module_defines_
