`timescale 1ns / 1ps
module key_schedule(
	input wire clk,
	input wire signal_start,
	output reg finished,
	input wire [127:0] key,
	input wire [63:0] round_ctr,
	output reg [127:0] outKey,
	output wire [3:0] state_response
    );
	 
	 
	 localparam widthshift_k0 = 3;
	 localparam widthshift_k1 = 8;
	 
	 localparam maxNrStates = 6;
	 parameter WAIT_FOR_START = 0;
	 parameter ASSIGNMENT = 1;
	 parameter SHIFT_k1 = 2;
	 parameter ADD_K0_K1 = 3;
	 parameter SHIFT_K0_XOR_P2 = 4;
	 parameter XOR_k1_k2 = 5;
	 parameter ASSIGN_RESULTS = 6;
	 
	 reg [3:0] state;
	 reg [63:0] k0;
	 reg [63:0] k1;
	 
	 localparam shiftwidth_p0 = 8;
	 localparam shiftwidth_p1 = 3;
	 	 
	 initial begin
		state <= 0;
		finished <= 0;
	end
	 
	 task inc_state;
	 begin
		if(state < maxNrStates) 
			state <= state + 1;
		else
			state <= 0;
	 end
	 endtask;
	 
	 function automatic [63:0] shift_right;
		 input [63:0] in;
		 input [4:0] shiftwidth;
		 begin
			shift_right = (in >>> shiftwidth) | (in <<< (64 - shiftwidth));
		 end
	 endfunction;
	 
	 function automatic [63:0] shift_left;
		 input [63:0] in;
		 input [4:0] shiftwidth;
		 begin
			shift_left = (in <<< shiftwidth) | (in >>> (64 - shiftwidth));
		 end
	 endfunction;
	 

	always @ (posedge clk) begin
		case (state)
			
			WAIT_FOR_START: begin
				if(signal_start)
					inc_state();
				finished <= 0;
			end
			
			ASSIGNMENT: begin
				k0 <= key[63:0];
				k1 <= key[127:64];
				inc_state();
			end
			
			SHIFT_k1: begin
				k0 <= shift_right(k0, 8);
				inc_state();
			end
			
			ADD_K0_K1: begin
				k0 <= k0 + k1;
				inc_state();
			end
			
			SHIFT_K0_XOR_P2: begin
				k1 <= shift_left(k1,3);
				k0 <= k0 ^ round_ctr;
				inc_state();
			end
			
			XOR_k1_k2: begin
				k1 <= k0 ^ k1;
				inc_state();
			end
			
			ASSIGN_RESULTS: begin
				outKey[63:0] <= k0;
				outKey[127:64] <= k1;
				inc_state();
				finished <= 1;
			end
			
		endcase;
		
	end
	
	assign state_response = state;




endmodule
