`ifndef _general_settings_
`define _general_settings_

	`define NR_ROUNDS 32'd31

`endif //_general_settings_
